module ROMControl (
    Addr,
    Data 
);
    parameter WIDTH_ADD = 6;
    parameter WIDTH_DATA = 20;
    input [WIDTH_ADD - 1:0] Addr;
    output reg [WIDTH_DATA - 1:0] Data;

    always @(Addr) begin
        case (Addr)
            //R type           
            6'd0:   Data = 20'b0_000_1_0_0_0_0000_0_00_000_01;
            6'd1:   Data = 20'b0_000_1_0_0_0_0001_0_00_000_01; 
            6'd2:   Data = 20'b0_000_1_0_0_0_0010_0_00_000_01;
            6'd3:   Data = 20'b0_000_1_0_0_0_0011_0_00_000_01;
            6'd4:   Data = 20'b0_000_1_0_0_0_0100_0_00_000_01; 
            6'd5:   Data = 20'b0_000_1_0_0_0_0101_0_00_000_01; 
            6'd6:   Data = 20'b0_000_1_0_0_0_0110_0_00_000_01; 
            6'd7:   Data = 20'b0_000_1_0_0_0_0111_0_00_000_01;
            6'd8:   Data = 20'b0_000_1_0_0_0_1000_0_00_000_01;
            6'd9:   Data = 20'b0_000_1_0_0_0_1001_0_00_000_01; 

            //I type
            6'd10:  Data = 20'b0_000_1_0_1_0_0000_0_00_000_01; 
            6'd11:  Data = 20'b0_000_1_0_1_0_0011_0_00_000_01; 
            6'd12:  Data = 20'b0_001_1_0_1_0_0100_0_00_000_01; 
            6'd13:  Data = 20'b0_000_1_0_1_0_0101_0_00_000_01;
            6'd14:  Data = 20'b0_000_1_0_1_0_1000_0_00_000_01; 
            6'd15:  Data = 20'b0_000_1_0_1_0_1001_0_00_000_01;  
            6'd16:  Data = 20'b0_010_1_0_1_0_0010_0_00_000_01; 
            6'd17:  Data = 20'b0_010_1_0_1_0_0110_0_00_000_01; 
            6'd18:  Data = 20'b0_010_1_0_1_0_0111_0_00_000_01; 

            //I type, Load Instruction
            6'd19:  Data = 20'b0_000_1_0_1_0_0000_0_00_000_00;
            6'd20:  Data = 20'b0_000_1_0_1_0_0000_0_00_001_00;
            6'd21:  Data = 20'b0_000_1_0_1_0_0000_0_00_010_00;
            6'd22:  Data = 20'b0_000_1_0_1_0_0000_0_00_011_00;
            6'd23:  Data = 20'b0_000_1_0_1_0_0000_0_00_100_00;

            //S type, Store Instruction
            6'd24:  Data = 20'b0_011_0_0_1_0_0000_1_00_000_00;
            6'd25:  Data = 20'b0_011_0_0_1_0_0000_1_01_000_00;
            6'd26:  Data = 20'b0_011_0_0_1_0_0000_1_11_000_00;

            //B type, Conditional Branch
            6'd27:  Data = 20'b1_100_0_0_1_1_0000_0_00_000_00;  //BEQ
            6'd28:  Data = 20'b0_100_0_0_1_1_0000_0_00_000_00;
            6'd29:  Data = 20'b0_100_0_0_1_1_0000_0_00_000_00;  //BNE
            6'd30:  Data = 20'b1_100_0_0_1_1_0000_0_00_000_00;
            6'd31:  Data = 20'b1_100_0_0_1_1_0000_0_00_000_00;  //BLT
            6'd32:  Data = 20'b0_100_0_0_1_1_0000_0_00_000_00;
            6'd33:  Data = 20'b0_100_0_0_1_1_0000_0_00_000_00;  //BGE
            6'd34:  Data = 20'b1_100_0_0_1_1_0000_0_00_000_00;
            6'd35:  Data = 20'b1_100_0_1_1_1_0000_0_00_000_00;  //BLTU
            6'd36:  Data = 20'b0_100_0_1_1_1_0000_0_00_000_00;
            6'd37:  Data = 20'b0_100_0_1_1_1_0000_0_00_000_00;  //BGEU
            6'd38:  Data = 20'b1_100_0_1_1_1_0000_0_00_000_00;

            //U type
            6'd39:  Data = 20'b0_101_1_0_1_0_1111_0_00_000_01;  //LUI
            6'd40:  Data = 20'b0_101_1_0_0_1_1110_0_00_000_01;  //AUIPC

            //J type, Unconditional Branch
            6'd41:  Data = 20'b1_110_1_0_1_1_0000_0_00_000_10;  //JAL
            6'd42:  Data = 20'b1_000_1_0_1_0_0000_0_00_000_10;  //JALR

            default: ;
        endcase
    end
endmodule